** sch_path: /ALL/git_olisnr/TO_Dec2024/RF_amplifiers/design_data/xschem/shunt_regulator/SHUNT_3V1.sch
**.subckt SHUNT_3V1 VSS VDD REFADJ REF1.2 SHUNT_GND
*.iopin VSS
*.iopin VDD
*.iopin REFADJ
*.iopin REF1.2
*.iopin SHUNT_GND
VDD net1 GND 5 ac 1
VSS GND VSS 0
Vzero 0 GND 0
Vmeas13 VDD net2 0
XM11 REF1.2 net8 net2 VDD sg13_hv_pmos w=8e-05 l=2e-06 ng=8
Vmeas14 net4 VSS 0
Vmeas15 net3 VSS 0
XQ3 net3 net3 net9 pnpMPA
XM12 net8 net7 net10 VSS sg13_hv_nmos w=1e-05 l=2e-06 ng=1
XM13 net7 net8 net5 VDD sg13_hv_pmos w=2e-05 l=2e-06 ng=2
XM14 net8 net8 net6 VDD sg13_hv_pmos w=2e-05 l=2e-06 ng=2
Vmeas16 VDD net5 0
Vmeas17 VDD net6 0
Vmeas18 net12 VSS 0
XM15 net7 net7 net12 VSS sg13_hv_nmos w=2e-06 l=2e-06 ng=1
XR9 net9 REF1.2 rppd w=1e-6 l=10e-6 m=1 b=10
XR10 net4 net10 rppd w=1e-6 l=10e-6 m=1 b=12
Vmeas7 net11 VSS 0
XM7 net17 net14 net11 VSS sg13_hv_nmos w=2e-06 l=2e-06 ng=1
Vmeas9 net13 VSS 0
XM6 net14 net14 net13 VSS sg13_hv_nmos w=2e-06 l=2e-06 ng=1
Vmeas10 VDD net15 0
XM8 net14 net8 net15 VDD sg13_hv_pmos w=2e-05 l=2e-06 ng=2
XM1 SHUNT_GND DRV_SHUNT net18 VDD sg13_hv_pmos w=0.0006 l=1e-06 ng=20
x12 net19 REF1.2 net16 VSS DRV_SHUNT net17 VDD DRV_SHUNT VDD VSS OTA3C nw=1e-06 nl=1e-06 pw=2e-06 pl=1e-06
XR1 net20 net16 rppd w=.5e-6 l=10e-6 m=1 b=14
XR2 net16 net21 rppd w=.5e-6 l=10e-6 m=1 b=10
Vmeas1 SHUNT_GND VSS 0
Vmeas2 net21 VSS 0
Vmeas3 VDD net20 0
Vmeas4 VDD net19 0
Vmeas5 VDD net18 0
XR3 REFADJ net10 rppd w=1e-6 l=10e-6 m=1 b=12
R4 VDD net1 100
XC4 REF1.2 VSS cap_cmim w=30.0e-6 l=30.0e-6
XC1 VDD net8 cap_cmim w=30.0e-6 l=30.0e-6
C2 VDD net22 1u
R5 net22 VSS 100m
**** begin user architecture code







* schematic: SHUNT_3V1
* dir:       /ALL/git_olisnr/TO_Dec2024/RF_amplifiers/design_data/xschem/shunt_regulator
* test:      /ALL/git_olisnr/TO_Dec2024/RF_amplifiers/design_data/xschem/shunt_regulator/OTA33_BiAS.sym

* mos_corner:
* mos_corner:






.option temp=27


.lib /home/ich/share/pdk/ihp-sg13g2/libs.tech/xyce/models/cornerRES.lib     res_typ
.lib /home/ich/share/pdk/ihp-sg13g2/libs.tech/xyce/models/cornerCAP.lib     cap_typ

.lib /home/ich/share/pdk/ihp-sg13g2/libs.tech/xyce/models/cornerMOShv.lib   mos_ss
.lib /home/ich/share/pdk/ihp-sg13g2/libs.tech/xyce/models/cornerMOSlv.lib   mos_ss
.lib /home/ich/share/pdk/ihp-sg13g2/libs.tech/xyce/models/cornerHBT.lib     hbt_typ

.param nw=1e-6
.param nl=1e-6
.param pw=2e-6
.param pl=1e-6
.param iset=3u

* .step dec iset 10u 100u 3

.dc temp -55 125 5
.print dc format=raw v(*) i(*)




**** end user architecture code
**.ends

* expanding   symbol:  /ALL/git_olisnr/TO_Dec2024/RF_amplifiers/design_data/xschem/shunt_regulator/OTA3C.sym # of pins=10
** sym_path: /ALL/git_olisnr/TO_Dec2024/RF_amplifiers/design_data/xschem/shunt_regulator/OTA3C.sym
** sch_path: /ALL/git_olisnr/TO_Dec2024/RF_amplifiers/design_data/xschem/shunt_regulator/OTA3C.sch
.subckt OTA3C VDD ip in VSS op sink C1 C3 C2 CGND  nw=1u nl=1u pw=2u pl=1u
*.ipin in
*.iopin VSS
*.iopin VDD
*.iopin sink
*.ipin ip
*.opin op
*.iopin C1
*.iopin C2
*.iopin C3
*.iopin CGND
XM1 net10 net18 net2 VDD sg13_hv_pmos w=2.4e-05 l=2e-06 ng=5 m=2
XM2 net9 net17 net2 VDD sg13_hv_pmos w=2.4e-05 l=2e-06 ng=5 m=2
Vmeas3 VDD net4 0
XM3 net10 net10 net1 VSS sg13_hv_nmos w=1e-06 l=1e-06 ng=1
XM4 net7 net10 net3 VSS sg13_hv_nmos w=2e-06 l=1e-06 ng=2
Vmeas8 net3 VSS 0
Vmeas9 net1 VSS 0
XM5 net8 V++ net4 VDD sg13_hv_pmos w=8e-06 l=1e-06 ng=2
**** begin user architecture code


**** end user architecture code
XM6 net2 V+ net8 VDD sg13_hv_pmos w=8e-06 l=1e-06 ng=2
XM7 net16 net9 net6 VSS sg13_hv_nmos w=2e-06 l=1e-06 ng=2
XM8 net9 net9 net5 VSS sg13_hv_nmos w=1e-06 l=1e-06 ng=1
Vmeas10 net5 VSS 0
Vmeas11 net6 VSS 0
XM9 net7 net17 net2 VDD sg13_hv_pmos w=2.4e-05 l=2e-06 ng=5 m=2
XM10 net16 net18 net2 VDD sg13_hv_pmos w=2.4e-05 l=2e-06 ng=5 m=2
Vmeas2 VDD net11 0
XM11 net14 net15 net11 VDD sg13_hv_pmos w=2e-06 l=1e-06 ng=1
XM12 op V+ net14 VDD sg13_hv_pmos w=2e-06 l=1e-06 ng=1
XM13 op V- net7 VSS sg13_hv_nmos w=1.5975e-05 l=1e-06 ng=9
Vmeas5 VDD net12 0
XM14 net13 net15 net12 VDD sg13_hv_pmos w=2e-06 l=1e-06 ng=1
XM15 net15 V+ net13 VDD sg13_hv_pmos w=2e-06 l=1e-06 ng=1
XM16 net15 V- net16 VSS sg13_hv_nmos w=1.5975e-05 l=1e-06 ng=9
x12 net19 sink V++ V+ V- V-- net20 OTA33_BiAS nw=1e-06 nl=1e-06 pw=2e-06 pl=1e-06
Vmeas1 net20 VSS 0
Vmeas4 VDD net19 0
R14 ip net18 1
R11 net17 in 1
XC2 C3 CGND cap_cmim w=9.0e-6 l=30.0e-6
XC3 C2 CGND cap_cmim w=9.0e-6 l=30.0e-6
XC4 C1 CGND cap_cmim w=9.0e-6 l=30.0e-6
.ends


* expanding   symbol:  /ALL/git_olisnr/TO_Dec2024/RF_amplifiers/design_data/xschem/shunt_regulator/OTA33_BiAS.sym # of pins=7
** sym_path: /ALL/git_olisnr/TO_Dec2024/RF_amplifiers/design_data/xschem/shunt_regulator/OTA33_BiAS.sym
** sch_path: /ALL/git_olisnr/TO_Dec2024/RF_amplifiers/design_data/xschem/shunt_regulator/OTA33_BiAS.sch
.subckt OTA33_BiAS VDD sink V++ V+ V- V-- VSS  nw=1u nl=1u pw=2u pl=1u
*.iopin VSS
*.iopin VDD
*.iopin sink
*.iopin V++
*.iopin V+
*.iopin V-
*.iopin V--
XM1 net4 V+ net2 VDD sg13_hv_pmos w=2e-06 l=1e-06 ng=2
Vmeas4 VDD net7 0
Vmeas6 net1 VSS 0
XM2 net3 V-- net1 VSS sg13_hv_nmos w=1e-06 l=1e-06 ng=1
XM3 V-- V- net3 VSS sg13_hv_nmos w=1e-06 l=1e-06 ng=1
XM4 net2 V++ net7 VDD sg13_hv_pmos w=2e-06 l=1e-06 ng=2
XM5 V- net4 V-- VSS sg13_hv_nmos w=1e-06 l=1e-06 ng=1
XM6 net4 net4 V- VSS sg13_hv_nmos w=1e-06 l=2e-06 ng=1
XM7 V++ V+ net5 VDD sg13_hv_pmos w=2e-06 l=1e-06 ng=2
XM8 net5 V++ net6 VDD sg13_hv_pmos w=2e-06 l=1e-06 ng=2
XM9 sink sink V+ VDD sg13_hv_pmos w=2e-06 l=2e-06 ng=1
XM10 V+ sink V++ VDD sg13_hv_pmos w=2e-06 l=1e-06 ng=2
Vmeas9 VDD net6 0
.ends

.GLOBAL GND
.end
